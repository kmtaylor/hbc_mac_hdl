#include <preprocessor/constants.vhh>

#ifndef RESET_BUTTON
#define RESET_BUTTON 0
#endif

#ifndef CLK_OUT
#define CLK_OUT 0
#endif

#ifndef USE_SWITCH
#define USE_SWITCH 0
#endif

#ifndef USE_8BIT_LED
#define USE_8BIT_LED 0
#endif

#ifndef USE_1BIT_LED
#define USE_1BIT_LED 0
#endif

#ifndef USE_LCD
#define USE_LCD 0
#endif

#ifndef USE_SPI
#define USE_SPI 0
#endif

#ifndef USE_BUTTON
#define USE_BUTTON 0
#endif

#ifndef USE_MEM
#define USE_MEM 0
#endif

#ifndef USE_MIG
#define USE_MIG 0
#endif

#ifndef USE_PAR_USB
#define USE_PAR_USB 0
#endif

#ifndef USE_FLASH
#define USE_FLASH 0
#endif

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library transceiver;
use transceiver.bits.all;

entity toplevel is
    port(
	clkin : in std_logic
#if RESET_BUTTON
	; rstbtn : in std_logic
#endif
	; s_data_out_filt : out std_logic
	; s_data_out_raw : out std_logic
	; s_data_in : in std_logic
#if CLK_OUT
	; serial_clk_out : out std_logic
#endif
#if USE_SWITCH
	; sw : in vec8_t
#endif
#if USE_8BIT_LED
	; Led : out vec8_t
#endif
#if USE_1BIT_LED
	; Led : out std_logic
#endif
#if USE_LCD
	; LCDD : inout vec8_t
	; LCDEN, LCDRW, LCDRS : out std_logic
#endif
#if USE_BUTTON
	; btn1, btn2 : in std_logic
#endif
#if USE_MEM
    #define MEM_DATA_WIDTH 16
    #define MEM_ADDR_WIDTH 13
    #define MEM_BYTES_WIDTH 2

	-- Physical memory interface
	; ddr2_dq	: inout std_logic_vector (MEM_DATA_WIDTH-1 downto 0)
	; ddr2_a	: out std_logic_vector (MEM_ADDR_WIDTH-1 downto 0)
	; ddr2_ba	: out std_logic_vector (1 downto 0)
	; ddr2_ras_n	: out std_logic
	; ddr2_cas_n	: out std_logic
	; ddr2_we_n	: out std_logic
	; ddr2_cs_n	: out std_logic
	; ddr2_cke	: out std_logic
	; ddr2_dm	: out std_logic_vector (MEM_BYTES_WIDTH-1 downto 0)
	; ddr2_dqs	: inout std_logic_vector (MEM_BYTES_WIDTH-1 downto 0)
#if USE_MIG
	; ddr2_odt	: out std_logic
	; ddr2_dqs_n	: inout std_logic_vector (MEM_BYTES_WIDTH-1 downto 0)
#endif
	; ddr2_ck	: out std_logic
	; ddr2_ck_n	: out std_logic
#endif
#if USE_PAR_USB
	-- USB Interface
	; UsbClk    : in std_logic
	; UsbEN	    : in std_logic
	; UsbEmpty  : in std_logic
	; UsbFull   : in std_logic
	; UsbOE	    : out std_logic
	; UsbAdr    : out std_logic_vector (1 downto 0)
	; UsbWR	    : out std_logic
	; UsbRD	    : out std_logic
	; UsbPktEnd : out std_logic
	; UsbDB	    : inout vec8_t
#endif
#if USE_SPI
	; hbc_ctrl_sclk : in std_logic
	; hbc_ctrl_mosi : in std_logic
	; hbc_ctrl_miso : out std_logic
	; hbc_data_sclk : in std_logic
	; hbc_data_mosi : in std_logic
	; hbc_data_miso : out std_logic
#endif
#if USE_PSOC
	; psoc_swdio : inout std_logic
	; psoc_swdck : inout std_logic
	; psoc_reset : inout std_logic
#endif
#if USE_FLASH
	; flash_sclk : out std_logic
	; flash_mosi : out std_logic
	; flash_miso : in std_logic
	; flash_ss : out std_logic
#endif
	);
end toplevel;

architecture toplevel_arch of toplevel is

    constant NUM_PERIPHERALS : natural := 9;
    constant PERIPH_HBC_TXFIFO	    : natural := 0;
    constant PERIPH_HBC_TXMOD	    : natural := 1;
    constant PERIPH_HBC_RXFIFO	    : natural := 2;
    constant PERIPH_HBC_SCRAMBLER   : natural := 3;
    constant PERIPH_MEM		    : natural := 4;
    constant PERIPH_SPI		    : natural := 5;
    constant PERIPH_FLASH_SPI	    : natural := 6;
    constant PERIPH_LCD		    : natural := 7;
    constant PERIPH_PAR_USB	    : natural := 8;

    type vec32n_t is array (NUM_PERIPHERALS-1 downto 0) of vec32_t;

    function peripheral_select (data : vec32n_t; ready : std_logic_vector) 
	return vec32_t is
    begin
	for i in ready'range loop
	    if ready(i) = '1' then
		return data(i);
	    end if;
	end loop;
	return (others => 'Z');
    end function peripheral_select;

    COMPONENT mcs_0
	PORT (
	    Clk : IN STD_LOGIC;
	    Reset : IN STD_LOGIC;
	    IO_Addr_Strobe : OUT STD_LOGIC;
	    IO_Read_Strobe : OUT STD_LOGIC;
	    IO_Write_Strobe : OUT STD_LOGIC;
	    IO_Address : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	    IO_Write_Data : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	    IO_Read_Data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	    IO_Ready : IN STD_LOGIC;
	    GPO1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
#if USE_8BIT_LED | USE_PSOC
	    GPO2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
#endif
	    GPI1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
#if USE_SWITCH | USE_PSOC
	    GPI2 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
#endif
	    INTC_Interrupt : IN STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
    END COMPONENT;
    
    constant RESET_DELAY : natural := 16;
#if !RESET_BUTTON
    signal rstbtn : std_logic;
#endif

    -- CPU interface
    signal io_read_strobe, io_write_strobe : std_logic;
    signal io_ready, io_addr_strobe : std_logic;
    signal io_address : vec32_t;
    signal io_write_data : vec32_t;
    signal io_read_data : vec32_t;
    signal irq_bus : std_logic_vector (15 downto 0);
    signal peripheral_data : vec32n_t;
    signal peripheral_ready : std_logic_vector (NUM_PERIPHERALS-1 downto 0);
    
    -- Internal memory signals
    signal phy_init_done    : std_logic;
    signal mem_fifo_full    : std_logic;
    signal rst0_tb	: std_logic;
    signal clk0_tb	: std_logic;
    signal app_wdf_afull    : std_logic;
    signal app_af_afull    : std_logic;
    signal rd_data_valid    : std_logic;
    signal app_rdf_rden    : std_logic;
    signal app_wdf_wren    : std_logic;
    signal app_af_wren    : std_logic;
    signal app_af_addr    : std_logic_vector (30 downto 0);
    signal app_af_cmd    : std_logic_vector (2 downto 0);
    signal rd_data_fifo_out    : std_logic_vector (127 downto 0);
    signal app_wdf_data    : std_logic_vector (127 downto 0);
    signal app_wdf_mask_data : std_logic_vector (15 downto 0);

    -- HBC data out mux
    signal s_data_out : std_logic;
    signal s_data_active : std_logic;
    signal s_data_out_switch : std_logic;
    
    -- HBC TX
    signal hbc_tx_fifo_flush : std_logic;
    signal hbc_tx_trigger : std_logic;
    signal hbc_tx_fifo_empty : std_logic;
    signal hbc_tx_fifo_almost_full : std_logic;
    signal hbc_tx_fifo_overflow : std_logic;

    -- HBC RX
    signal hbc_rx_fifo_almost_full : std_logic;
    signal hbc_rx_fifo_empty : std_logic;
    signal hbc_rx_enable : std_logic;
    signal hbc_rx_active : std_logic;
    signal hbc_rx_pkt_ready : std_logic;
    signal hbc_rx_pkt_ack : std_logic;

    -- PAR_USB
    signal usb_pkt_end : std_logic;
    signal usb_irq : std_logic;
    signal usb_clk : std_logic;
    
    -- Scrambler
    signal scram_reseed, scram_seed_val, scram_seed_clk : std_logic;

    -- Infrastructure
    signal serial_reset : std_logic;
    signal cpu_reset : std_logic;
    signal c_reset_shift_r : std_logic_vector(RESET_DELAY-1 downto 0);
    signal s_reset_shift_r : std_logic_vector(RESET_DELAY-1 downto 0);
    attribute equivalent_register_removal : string;
    attribute max_fanout : string;
    attribute shreg_extract : string;
    attribute equivalent_register_removal of cpu_reset : signal is "no";
    attribute max_fanout of cpu_reset : signal is "10";
    attribute shreg_extract of cpu_reset : signal is "no";
    attribute equivalent_register_removal of serial_reset : signal is "no";
    attribute max_fanout of serial_reset : signal is "10";
    attribute shreg_extract of serial_reset : signal is "no";
    signal clk_debounce, clkin_ibufg : std_logic;
    signal pll_clk, cpu_clk, serial_clk, serial_clk_90 : std_logic;
    signal serial_clk_tmp : std_logic;
    signal mem_clk0, mem_clk90, mem_clkdiv0, mem_clk200 : std_logic;
    signal pll_locked, mem_pll_locked : std_logic;
    signal serial_dcm_locked : std_logic;
    signal cpu_dcm_locked : std_logic;
    signal clk_lock_int : std_logic;

    -- PSOC HSSP interface
    signal psoc_swdio_dir, psoc_swdck_dir, psoc_xres_dir : std_logic;
    signal psoc_swdio_i, psoc_swdck_i, psoc_xres_i : std_logic;
    signal psoc_swdio_o, psoc_swdck_o, psoc_xres_o : std_logic;

    -- SPI interface
    signal hbc_ctrl_spi_int, hbc_data_spi_int : std_logic;

    signal btn1_d : std_logic;
    signal btn2_d : std_logic;

begin

#if !RESET_BUTTON
    rstbtn <= '1';
#endif
    
    cpu_reset_sync_proc : process (cpu_clk, rstbtn) begin
        if rstbtn = '0' then
            c_reset_shift_r <= (others => '1');
        elsif cpu_clk'event and cpu_clk = '1' then
	    c_reset_shift_r <= shift_left(c_reset_shift_r, 1);
        end if;
    end process cpu_reset_sync_proc;

    cpu_reset <= c_reset_shift_r(RESET_DELAY-1);

    serial_reset_sync_proc : process (serial_clk, rstbtn) begin
        if rstbtn = '0' then
            s_reset_shift_r <= (others => '1');
        elsif serial_clk'event and serial_clk = '1' then
	    s_reset_shift_r <= shift_left(s_reset_shift_r, 1);
        end if;
    end process serial_reset_sync_proc;

    serial_reset <= s_reset_shift_r(RESET_DELAY-1);

#if CLK_OUT
    serial_clk_out <= serial_clk;
#endif

    cpu_clk <= mem_clk0;

    clk_lock_int <= not(pll_locked and serial_dcm_locked and 
		cpu_dcm_locked and mem_pll_locked);

#if USE_MIG
    mem_fifo_full <= app_af_afull or app_wdf_afull;
#else
    mem_fifo_full <= '0';
#endif

#if XILINX_VIRTEX
    -- 100MHz XTal to 42MHz PLL
    core_pll : entity work.pll_core
	port map (
	    CLKIN1_IN => clkin,
	    RST_IN => '0',
	    CLKOUT0_OUT => pll_clk,
	    CLKIN_IBUFG => clkin_ibufg,
	    LOCKED_OUT => pll_locked);

    -- 100MHz XTal to 125MHz Mem clock (Also 200MHz and 62.5MHz)
    mem_pll : entity work.pll_mem
	port map (
	    CLKIN1_IN => clkin_ibufg,
	    RST_IN => '0',
	    CLKOUT0_OUT => mem_clk0,
	    CLKOUT1_OUT => mem_clk90,
	    CLKOUT2_OUT => mem_clkdiv0,
	    CLKOUT3_OUT => mem_clk200,
	    LOCKED_OUT => mem_pll_locked);

#if USE_PAR_USB
    usb_bufr : component BUFR
	port map (
	    I => UsbClk,
	    O => usb_clk);
#endif
    
    cpu_dcm_locked <= '1';

#define SERIAL_DIV 0
#if SERIAL_DIV
    clk_div_1 : entity work.clock_divider
	generic map (DIV_BY => 8)
	port map (clk => serial_clk_tmp, clk_div => serial_clk);

    -- 42MHz PLL to 42MHz serial clock for TX
    serial_clk_dcm : entity work.dcm_serial
	port map (
	    CLKIN_IN => pll_clk,
	    RST_IN => '0',
	    CLK0_OUT => serial_clk_tmp,
	    CLK90_OUT => serial_clk_90,
	    LOCKED_OUT => serial_dcm_locked);
#else
    -- 42MHz PLL to 42MHz serial clock for TX
    serial_clk_dcm : entity work.dcm_serial
	port map (
	    CLKIN_IN => pll_clk,
	    RST_IN => '0',
	    CLK0_OUT => serial_clk,
	    CLK90_OUT => serial_clk_90,
	    LOCKED_OUT => serial_dcm_locked);
#endif
#endif /* -- XILINX_VIRTEX */

#if XILINX_SPARTAN
    -- 62.5MHz XTal to 100MHz PLL
    mem_pll : entity work.pll_mem
	port map (
	    CLKIN1_IN => clkin,
	    RST_IN => '0',
	    CLKOUT0_OUT => mem_clk0,
	    CLKOUT1_OUT => mem_clk90,
	    LOCKED_OUT => pll_locked);

    mem_pll_locked <= '1';
    cpu_dcm_locked <= '1';

    -- 100MHz to 42MHz PLL serial clock for TX
    serial_clk_pll : entity work.pll_serial
	port map (
	    CLKIN1_IN => mem_clk0,
	    RST_IN => '0',
	    CLKOUT0_OUT => serial_clk,
	    CLKOUT1_OUT => serial_clk_90,
	    LOCKED_OUT => serial_dcm_locked);
#endif /* -- XILINX_SPARTAN */
	    
#if USE_BUTTON
    -- 125MHz cpu_clk to 6.25kHz clk for pushbutton debouncing 
    clk_div_0 : entity work.clock_divider
	generic map (DIV_BY => 20E3)
	port map (clk => cpu_clk, clk_div => clk_debounce);
#endif
	    
    cpu_0 : component mcs_0
	port map (
	    Clk => cpu_clk,
	    Reset => cpu_reset,
	    IO_Addr_Strobe => io_addr_strobe,
	    IO_Read_Strobe => io_read_strobe,
	    IO_Write_Strobe => io_write_strobe,
	    IO_Address => io_address,
	    IO_Write_Data => io_write_data,
	    IO_Read_Data => io_read_data,
	    IO_Ready => io_ready,
#if USE_SWITCH
	    GPI2 => sw,
#endif
	    GPO(HBC_TX_TRIGGER, hbc_tx_trigger),
	    GPO(HBC_TX_FLUSH, hbc_tx_fifo_flush),
	    GPO(SCRAM_RESEED, scram_reseed),
	    GPO(SCRAM_SEED_VAL, scram_seed_val),
	    GPO(SCRAM_SEED_CLK, scram_seed_clk),
	    GPO(HBC_RX_PKT_ACK, hbc_rx_pkt_ack),
	    GPO(HBC_RX_ENABLE, hbc_rx_enable),
#if USE_1BIT_LED
	    GPO(LED_1BIT, led),
#elif USE_PAR_USB
	    GPO(USB_PKT_END, usb_pkt_end),
#else
	    GPO1(7) => open,
#endif
#if USE_8BIT_LED
	    GPO2 => Led,
#endif
#if USE_PSOC
	    GPI(PSOC_DATA, psoc_swdio_i),
	    GPI(PSOC_CLOCK, psoc_swdck_i),
	    GPI(PSOC_RESET, psoc_xres_i),
	    GPI2(7 downto 3) => (others => '0'),
	    GPO(PSOC_DATA, psoc_swdio_o),
	    GPO(PSOC_DATA_DIR, psoc_swdio_dir),
	    GPO(PSOC_CLOCK, psoc_swdck_o),
	    GPO(PSOC_CLOCK_DIR, psoc_swdck_dir),
	    GPO(PSOC_RESET, psoc_xres_o),
	    GPO(PSOC_RESET_DIR, psoc_xres_dir),
#else
	    GPO2(5 downto 0) => open,
#endif
#if USE_FLASH
	    GPO(FLASH_SS, flash_ss),
#else
	    GPO2(6) => open,
#endif
	    GPO(HBC_DATA_SWITCH, s_data_out_switch),
	    INTC_Interrupt => irq_bus,
	    GPI1 => irq_bus);

    IRQ(IRQ_BUTTON, btn1_d);
    IRQ(IRQ_TX_FIFO_EMPTY, hbc_tx_fifo_empty);
    IRQ(IRQ_TX_FIFO_ALMOST_FULL, hbc_tx_fifo_almost_full);
    IRQ(IRQ_TX_FIFO_OVERFLOW, hbc_tx_fifo_overflow);
    IRQ(IRQ_RX_ACTIVE, hbc_rx_active);
    IRQ(IRQ_RX_DATA_READY, not(hbc_rx_fifo_empty));
    IRQ(IRQ_RX_PKT_READY, hbc_rx_pkt_ready);
    IRQ(IRQ_RX_FIFO_ALMOST_FULL, hbc_rx_fifo_almost_full);
    IRQ(IRQ_CLOCK_LOSS, clk_lock_int);
    IRQ(IRQ_RAM_INIT, not(phy_init_done));
    IRQ(IRQ_RAM_FIFO_FULL, mem_fifo_full);
    IRQ(IRQ_BUTTON_2, btn2_d);
#if USE_PAR_USB
    IRQ(IRQ_USB_INT, usb_irq);
    IRQ(IRQ_USB_FULL, UsbFull);
    IRQ(IRQ_USB_EN, UsbEN);
    IRQ(IRQ_USB_EMPTY, UsbEmpty);
#elif USE_SPI
    IRQ(IRQ_HBC_CTRL_SPI, hbc_ctrl_spi_int);
    IRQ(IRQ_HBC_DATA_SPI, hbc_data_spi_int);
#endif

    io_read_data <= peripheral_select(peripheral_data, peripheral_ready);
    io_ready <= bool_to_bit(peripheral_ready /= zeros(peripheral_ready'length));
    
    mem_if : entity work.mem_interface
	port map (
	    cpu_clk => cpu_clk,
	    reset => cpu_reset,
	    io_addr => io_address (7 downto 0),
	    io_d_in => io_write_data,
	    io_d_out => peripheral_data(PERIPH_MEM),
	    io_addr_strobe => io_addr_strobe,
	    io_read_strobe => io_read_strobe,
	    io_write_strobe => io_write_strobe,
	    io_ready => peripheral_ready(PERIPH_MEM),
	    app_af_cmd => app_af_cmd,
	    app_af_addr => app_af_addr,
	    app_af_wren => app_af_wren,
	    app_wdf_data => app_wdf_data,
	    app_wdf_wren => app_wdf_wren,
	    app_wdf_mask_data => app_wdf_mask_data,
	    rd_data_valid => rd_data_valid,
	    rd_data_fifo_out => rd_data_fifo_out);
	    
#if USE_MIG
    ram : entity work.mem_controller
	port map (
	    -- Physical RAM interface
	    ddr2_dq		=> ddr2_dq,
	    ddr2_a		=> ddr2_a,
	    ddr2_ba		=> ddr2_ba,
	    ddr2_ras_n		=> ddr2_ras_n,
	    ddr2_cas_n		=> ddr2_cas_n,
	    ddr2_we_n		=> ddr2_we_n,
	    ddr2_cs_n		=> ddr2_cs_n,
	    ddr2_odt		=> ddr2_odt,
	    ddr2_cke		=> ddr2_cke,
	    ddr2_dm		=> ddr2_dm,
	    ddr2_dqs		=> ddr2_dqs,
	    ddr2_dqs_n		=> ddr2_dqs_n,
	    ddr2_ck		=> ddr2_ck,
	    ddr2_ck_n		=> ddr2_ck_n,
	    -- Infrastructure
	    clk0		=> mem_clk0,
	    clk90		=> mem_clk90,
	    clkdiv0		=> mem_clkdiv0,
	    clk200		=> mem_clk200,
	    locked		=> mem_pll_locked,
	    sys_rst_n		=> rstbtn,
	    phy_init_done	=> phy_init_done,
	    rst0_tb		=> rst0_tb,
	    clk0_tb		=> clk0_tb,
	    -- Address FIFO
	    app_af_cmd		=> app_af_cmd,
	    app_af_addr		=> app_af_addr,
	    app_af_wren		=> app_af_wren,
	    app_af_afull	=> app_af_afull,
	    -- Write FIFO
	    app_wdf_data	=> app_wdf_data,
	    app_wdf_wren	=> app_wdf_wren,
	    app_wdf_afull	=> app_wdf_afull,
	    app_wdf_mask_data	=> app_wdf_mask_data,
	    --Read FIFO
	    rd_data_valid	=> rd_data_valid,
	    rd_data_fifo_out	=> rd_data_fifo_out);
#endif

#if USE_MEM
    ram : entity work.ddr
	port map (
	    mem_clk => mem_clk0,
	    reset_i => cpu_reset,
	    app_af_cmd => app_af_cmd(0),
	    app_af_addr(30 downto 0) => app_af_addr,
	    app_af_addr(31) => '0',
	    app_wdf_data => app_wdf_data(31 downto 0),
	    app_af_wren => app_af_wren,
	    app_wdf_mask_data => app_wdf_mask_data(3 downto 0),
	    rd_data_valid => rd_data_valid,
	    rd_data_fifo_out => rd_data_fifo_out(31 downto 0),

	    ram_clk => ddr2_ck,
	    ram_clk_n => ddr2_ck_n,
	    ram_cke => ddr2_cke,
	    ram_cs_n => ddr2_cs_n,
	    ram_cmd(0) => ddr2_we_n,
	    ram_cmd(1) => ddr2_cas_n,
	    ram_cmd(2) => ddr2_ras_n,
	    ram_ba => ddr2_ba,
	    ram_addr => ddr2_a,
	    ram_dm => ddr2_dm,
	    ram_dqs => ddr2_dqs,
	    ram_dq => ddr2_dq);

    phy_init_done <= '1';
#endif

    hbc_tx: entity work.hbc_tx
	port map (
	    cpu_clk => cpu_clk,
	    cpu_reset => cpu_reset,
	    serial_clk => serial_clk,
	    serial_reset => serial_reset,
	    io_addr => io_address (7 downto 0),
	    io_d_in => io_write_data,
	    io_d_out => peripheral_data(PERIPH_HBC_TXFIFO),
	    io_addr_strobe => io_addr_strobe,
	    io_read_strobe => io_read_strobe,
	    io_write_strobe => io_write_strobe,
	    io_ready_fifo => peripheral_ready(PERIPH_HBC_TXFIFO),
	    io_ready_mod => peripheral_ready(PERIPH_HBC_TXMOD),
	    hbc_tx_fifo_flush => hbc_tx_fifo_flush,
	    hbc_tx_trigger => hbc_tx_trigger,
	    hbc_tx_fifo_empty => hbc_tx_fifo_empty,
	    hbc_tx_fifo_almost_full => hbc_tx_fifo_almost_full,
	    hbc_tx_fifo_overflow => hbc_tx_fifo_overflow,
	    s_data_active => s_data_active,
	    s_data_out => s_data_out);

    s_data_out_mux : process (s_data_out_switch,
				     s_data_out, s_data_active) begin
	if s_data_out_switch = '1' then
	    s_data_out_filt <= 'Z';
	    if s_data_active = '1' then
		s_data_out_raw <= s_data_out;
	    else
		s_data_out_raw <= 'Z';
	    end if;
	else
	    if s_data_active = '1' then
		s_data_out_filt <= s_data_out;
	    else
		s_data_out_filt <= 'Z';
	    end if;
	    s_data_out_raw <= 'Z';
	end if;
    end process s_data_out_mux;

    hbc_rx: entity work.hbc_rx
	port map (
	    cpu_clk => cpu_clk,
	    cpu_reset => cpu_reset,
	    serial_clk => serial_clk,
	    serial_clk_90 => serial_clk_90,
	    serial_reset => serial_reset,
	    io_addr => io_address (7 downto 0),
	    io_d_out => peripheral_data(PERIPH_HBC_RXFIFO),
	    io_addr_strobe => io_addr_strobe,
	    io_read_strobe => io_read_strobe,
	    io_ready => peripheral_ready(PERIPH_HBC_RXFIFO),
	    hbc_rx_enable => hbc_rx_enable,
	    hbc_rx_active => hbc_rx_active,
	    hbc_rx_fifo_almost_full => hbc_rx_fifo_almost_full,
	    hbc_rx_fifo_empty => hbc_rx_fifo_empty,
	    hbc_rx_pkt_ready => hbc_rx_pkt_ready,
	    hbc_rx_pkt_ack => hbc_rx_pkt_ack,
	    s_data_in => s_data_in);

    scrambler : entity work.scrambler
	port map (
	    cpu_clk => cpu_clk,
	    reset => cpu_reset,
	    reseed => scram_reseed,
	    seed_val => scram_seed_val,
	    seed_clk => scram_seed_clk,
	    io_addr => io_address (7 downto 0),
	    io_d_out => peripheral_data(PERIPH_HBC_SCRAMBLER),
	    io_addr_strobe => io_addr_strobe,
	    io_read_strobe => io_read_strobe,
	    io_ready => peripheral_ready(PERIPH_HBC_SCRAMBLER));

#if USE_SPI
    spi_hbc : entity work.spi_interface
	port map (
	    clk => cpu_clk,
	    reset => cpu_reset,
	    io_addr => io_address (7 downto 0),
	    io_d_out => peripheral_data(PERIPH_SPI),
	    io_d_in => io_write_data,
	    io_addr_strobe => io_addr_strobe,
	    io_read_strobe => io_read_strobe,
	    io_write_strobe => io_write_strobe,
	    io_ready => peripheral_ready(PERIPH_SPI),
	    hbc_data_int => hbc_data_spi_int,
	    hbc_ctrl_int => hbc_ctrl_spi_int,
	    hbc_data_sclk => hbc_data_sclk,
	    hbc_data_mosi => hbc_data_mosi,
	    hbc_data_miso => hbc_data_miso,
	    hbc_data_ss => psoc_swdck,
	    hbc_ctrl_sclk => hbc_ctrl_sclk,
	    hbc_ctrl_mosi => hbc_ctrl_mosi,
	    hbc_ctrl_miso => hbc_ctrl_miso,
	    hbc_ctrl_ss => psoc_swdio);
#endif

#if USE_PSOC
    psoc_interface : entity work.psoc_interface
	port map (
	    swdio_dir => psoc_swdio_dir,
	    swdck_dir => psoc_swdck_dir,
	    xres_dir => psoc_xres_dir,
	    swdio_i => psoc_swdio_i,
	    swdio_o => psoc_swdio_o,
	    swdck_i => psoc_swdck_i,
	    swdck_o => psoc_swdck_o,
	    xres_i => psoc_xres_i,
	    xres_o => psoc_xres_o,
	    swdio => psoc_swdio,
	    swdck => psoc_swdck,
	    xres => psoc_reset);
#endif

#if USE_FLASH
    flash_interface : entity work.flash_interface
	generic map (DIVIDER => 10)
	port map (
	    cpu_clk => cpu_clk,
	    reset => cpu_reset,
	    io_addr => io_address (7 downto 0),
	    io_d_in => io_write_data,
	    io_d_out => peripheral_data(PERIPH_FLASH_SPI),
	    io_addr_strobe => io_addr_strobe,
	    io_read_strobe => io_read_strobe,
	    io_write_strobe => io_write_strobe,
	    io_ready => peripheral_ready(PERIPH_FLASH_SPI),
	    flash_sclk => flash_sclk,
	    flash_mosi => flash_mosi,
	    flash_miso => flash_miso,
	    flash_ss => open);
#endif

#if USE_PAR_USB
    usb_0 : entity work.usb_fifo
	port map (
	    usb_clk => usb_clk,
	    cpu_clk => cpu_clk,
	    reset => cpu_reset,
	    io_addr => io_address (7 downto 0),
	    io_d_in => io_write_data,
	    io_d_out => peripheral_data(PERIPH_PAR_USB),
	    io_addr_strobe => io_addr_strobe,
	    io_read_strobe => io_read_strobe,
	    io_write_strobe => io_write_strobe,
	    io_ready => peripheral_ready(PERIPH_PAR_USB),
	    pkt_end => usb_pkt_end,
	    UsbIRQ => usb_irq,
	    UsbDB => UsbDB,
	    UsbAdr => UsbAdr,
	    UsbOE => UsbOE,
	    UsbWR => UsbWR,
	    UsbRD => UsbRD,
	    UsbPktEnd => UsbPktEnd,
	    UsbEmpty => UsbEmpty,
	    UsbFull => UsbFull,
	    UsbEN => UsbEN,
	    UsbDBG => open);
#endif

#if USE_LCD
    lcd_0 : entity work.lcd_interface
	port map (
	    clk => cpu_clk,
	    reset => cpu_reset,
	    io_addr => io_address (7 downto 0),
	    io_d_in => io_write_data,
	    io_d_out => peripheral_data(PERIPH_LCD),
	    io_addr_strobe => io_addr_strobe,
	    io_read_strobe => io_read_strobe,
	    io_write_strobe => io_write_strobe,
	    io_ready => peripheral_ready(PERIPH_LCD),
	    lcd_data => LCDD,
	    lcd_en => LCDEN,
	    lcd_rw => LCDRW,
	    lcd_rs => LCDRS);
#endif
	
#if USE_BUTTON
    db_btn1 : entity work.debounce
	port map (
	    clk => clk_debounce,
	    d_in => btn1,
	    q_out => btn1_d);

    db_btn2 : entity work.debounce
	port map (
	    clk => clk_debounce,
	    d_in => btn2,
	    q_out => btn2_d);
#else
    btn1_d <= '0';
    btn2_d <= '0';
#endif

end toplevel_arch;

