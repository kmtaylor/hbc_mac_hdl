#include <preprocessor/constants.vhh>
#include "send_packet.vhh"

#ifndef STIMULUS
#define STIMULUS 1
#endif

#ifndef SERIAL_CLK_NS
#define SERIAL_CLK_NS 23.81
#endif

library ieee;
use ieee.std_logic_1164.all;

entity transmitter_tb is
#if !STIMULUS
    port (
	clk, serial_clk, reset, parallel_to_serial_enable : in std_logic;
	fi_write_strobe, fi_addr_strobe : in std_logic;
	fi_d : in std_logic_vector (31 downto 0);
	fi_addr : in std_logic_vector (7 downto 0);
	io_write_strobe, io_addr_strobe : in std_logic;
	io_d_in : in std_logic_vector (31 downto 0);
	io_addr : in std_logic_vector (7 downto 0);
	io_ready : out std_logic;
	prog_full : out std_logic;
	s_data_out : out std_logic);
#endif
end transmitter_tb;
 
architecture testbench of transmitter_tb is 
 
    component fifo_tx port (
        rst : IN STD_LOGIC;
        wr_clk : IN STD_LOGIC;
        rd_clk : IN STD_LOGIC;
        din : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        wr_en : IN STD_LOGIC;
        rd_en : IN STD_LOGIC;
        dout : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        full : OUT STD_LOGIC;
	prog_full : OUT STD_LOGIC;
        overflow : OUT STD_LOGIC;
        empty : OUT STD_LOGIC;
        underflow : OUT STD_LOGIC);
    end component fifo_tx;

   --Inputs
#if STIMULUS
    signal clk : std_logic := '0';
    signal reset : std_logic := '0';
    signal io_addr : std_logic_vector(7 downto 0) := (others => '0');
    signal io_d_in : std_logic_vector(31 downto 0) := (others => '0');
    signal io_addr_strobe : std_logic := '0';
    signal io_write_strobe : std_logic := '0';
    signal io_ready : std_logic;
#endif
    signal io_read_strobe : std_logic := '0';
    signal sub_io_ready : std_logic;

    signal tmp_addr : std_logic_vector (7 downto 0);
    signal tmp_d : std_logic_vector (31 downto 0);
    signal tmp_addr_strobe : std_logic;
    signal tmp_write_strobe : std_logic;

#if STIMULUS
    signal fi_addr : std_logic_vector (7 downto 0) := (others => '0');
    signal fi_d : std_logic_vector (31 downto 0) := (others => '0');
    signal fi_addr_strobe : std_logic := '0';
    signal fi_write_strobe : std_logic := '0';
#endif

    --Outputs
    signal sub_addr_out: std_logic_vector (7 downto 0);
    signal sub_d_out   : std_logic_vector (31 downto 0);
    signal sub_addr_strobe : std_logic;
    signal sub_write_strobe : std_logic;
    signal bus_master : std_logic;

    signal cho_demod_out : std_logic;

    -- FIFO
    signal fifo_d_out : std_logic_vector (31 downto 0);
    signal fifo_wren, fifo_rden : std_logic;
    signal full, overflow, empty, underflow : std_logic;
    signal from_fifo : std_logic_vector (31 downto 0);
#if STIMULUS
    signal prog_full : std_logic;
#endif

    -- P2S
#if STIMULUS
    signal serial_clk, parallel_to_serial_enable : std_logic;
    signal s_data_out : std_logic;
#endif

    -- Clock period definitions
    constant clk_period : time := 10 ns;
    constant s_clk_period : time := SERIAL_CLK_NS ns;
    
#if STIMULUS
    type val_ft is file of std_logic;
    type time_ft is file of time;
    file val_file : val_ft open WRITE_MODE is "tx_data.value";
    file time_file : time_ft open WRITE_MODE is "tx_data.time";
    procedure write_val(val : std_logic) is begin
        write(val_file, val);
        write(time_file, now);
    end procedure write_val;
#endif
begin
 
    cho_demod : entity work.cho_demod port map (
	clk => serial_clk,
	data => s_data_out,
	output => cho_demod_out);

    -- Instantiate the Unit Under Test (UUT)
    modulator : entity work.modulator port map (
	clk => clk,
	reset => reset,
	io_addr => io_addr,
	io_d_in => io_d_in,
	io_addr_strobe => io_addr_strobe,
	io_write_strobe => io_write_strobe,
	io_ready => io_ready,
	bus_master => bus_master,
	sub_addr_out => sub_addr_out,
	sub_d_out => sub_d_out,
	sub_addr_strobe => sub_addr_strobe,
	sub_write_strobe => sub_write_strobe,
	sub_io_ready => sub_io_ready,
	fifo_almost_full => prog_full);

    process (bus_master, sub_addr_out, sub_d_out, sub_addr_strobe,
		    sub_write_strobe, fi_addr, fi_d, fi_addr_strobe,
		    fi_write_strobe) begin
	if bus_master = '1' then
	    tmp_addr <= sub_addr_out;
	    tmp_d <= sub_d_out;
	    tmp_addr_strobe <= sub_addr_strobe;
	    tmp_write_strobe <= sub_write_strobe;
	else
	    tmp_addr <= fi_addr;
	    tmp_d <= fi_d;
	    tmp_addr_strobe <= fi_addr_strobe;
	    tmp_write_strobe <= fi_write_strobe;
	end if;
    end process;

    tx_fifo_interface : entity work.tx_fifo_interface port map (
	clk => clk,
	reset => reset,
	trigger => '0',
	io_addr => tmp_addr,
	io_d_in => tmp_d,
	io_d_out => open,
	io_addr_strobe => tmp_addr_strobe,
	io_read_strobe => '0',
	io_write_strobe => tmp_write_strobe,
	io_ready => sub_io_ready,
	fifo_d_out => fifo_d_out,
	fifo_d_in => (others => '0'),
	fifo_wren => fifo_wren,
	fifo_rden => open);

    p_to_s : entity work.parallel_to_serial port map (
	clk => serial_clk,
	reset => reset,
	trigger => parallel_to_serial_enable,
	trig_clk => clk,
	fifo_d_in => from_fifo,
	fifo_rden => fifo_rden,
	fifo_empty => empty,
	data_out => s_data_out);

    tx_fifo : component fifo_tx port map (
        rst => reset,
        wr_clk => clk,
        rd_clk => serial_clk,
        din => fifo_d_out,
        wr_en => fifo_wren,
        rd_en => fifo_rden,
        dout => from_fifo,
        full => full,
	prog_full => prog_full,
        overflow => overflow,
        empty => empty,
        underflow => underflow);

#if STIMULUS
    -- Clock process definitions
    clk_process : process begin
	clk <= '0';
	wait for clk_period/2;
	clk <= '1';
	wait for clk_period/2;
    end process;

    s_clk_process : process begin
	serial_clk <= '0';
	wait for s_clk_period/2;
	serial_clk <= '1';
	wait for s_clk_period/2;
    end process;
#endif

#if STIMULUS
    -- Stimulus process
    stim_proc: process begin	
	-- hold reset state for 60 ns.
	reset <= '1';
	parallel_to_serial_enable <= '0';
	wait for 60 ns;
	reset <= '0';

	wait for clk_period * 5.5;

	-- Trigger P2S
	TRIGGER()
	SEND_PACKET()

	wait;
    end process;
#endif

#if STIMULUS
    write_proc : process(s_data_out) begin
	write_val(s_data_out);
    end process;
#endif

end;
